module IMEM (
    input [31:0] addr,
    output [31:0] inst
);
    reg [31:0] memory [0:255];
    
    assign inst = memory[addr[31:2]];

    always @(*) begin
        $display("IMEM: Cycle=%0d, addr=%h, inst=%h", $time/10, addr, inst);
    end
endmodule